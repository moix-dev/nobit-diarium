module main

fn test_main() {
    assert true
}